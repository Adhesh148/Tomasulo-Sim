`include "fpMult.v"

module top;
	reg[31:0] X1,X2;
	wire[31:0] X3;

	fpMult fp_0 (X3 ,X1, X2);

	// Setup the monitoring for the signal values
	initial
	begin
		$monitor($time," X1 = %b,  X2 = %b --- X3 = %b\n",X1,X2,X3);
		$dumpfile("fpM.vcd");
		$dumpvars;
	end

	// Simulate the inputs
	initial
	begin
		X1 = 0; X2 = 0;

		// 9.75 * 0.5625 = 5.484375
		#5 X2 = 32'b01000001000111000000000000000000; X1 = 32'b00111111000100000000000000000000;

		// 4 * 0.10000000149 = 0.40000000596
		#5 X2 = 32'b01000000100000000000000000000000; X1 = 32'b00111101110011001100110011001101;

		// 4 * -0.25 = -1 
		#5 X1 = 32'b01000000100000000000000000000000; X2 = 32'b10111110100000000000000000000000;

		// 4.13000011444 * 2.40000009537 = 9.91200065613
		#5 X1 = 32'b01000000100001000010100011110110; X2 = 32'b01000000000110011001100110011010;

		// -4.0 * 0.25 = -1
		#5 X1 = 32'b11000000100000000000000000000000; X2 = 32'b00111110100000000000000000000000;

		// 4 * -6.25 = -25
		#5 X1 = 32'b01000000100000000000000000000000; X2 = 32'b11000000110010000000000000000000;

		// 4 * -4 = -16.0
		#5 X1 = 32'b01000000100000000000000000000000; X2 = 32'b11000000100000000000000000000000;

		// -4 * (-4.0078125) = 16.03125
		#5 X1 = 32'b11000000100000000000000000000000; X2 = 32'b11000000100000000100000000000000;

		// -2312.12 * (-142.912) = 330429.6875
		#5 X1 = 32'b11000101000100001000000111101100; X2 = 32'b11000011000011101110100101111001;
		
		// -990.99 * 0.99 = -981.080078125
		#5 X1 = 32'b11000100011101111011111101011100; X2 = 32'b00111111011111010111000010100100;

		// -6.13802377216e+11 * -1.53450594304e+11 = 9.418833665e+22
		#5 X1 = 32'b11010011000011101110100101111001; X2 = 32'b11010010000011101110100101111001;

		// 0 * x = 0
		#5 X1 = 32'b00000000000000000000000000000000; X2 = 32'b11010010000011101110100101111001;

		//  nan * 0 = nan
		#5 X1 = 32'b01111111111111111111111111111111; X2 = 32'b00000000000000000000000000000000;

		//  inf * 0 = nan
		#5 X1 = 32'b01111111100000000000000000000000; X2 = 32'b00000000000000000000000000000000;

		//  nan * inf = nan
		#5 X1 = 32'b01111111111111111111111111111111; X2 = 32'b01111111100000000000000000000000;
	end

endmodule