module parallelPrefixCkt(Y,A,B);
	output reg[1:0] Y;
	input[1:0] A,B;

	always @(A or B)
	begin
		if(A == 2'b00 || A == 2'b11)
			assign Y = A;
		else
			assign Y = B;
	end
endmodule

module doublingCLA_64(Sum,Cout,A,B,Cin);

	// I/O Port Declarations
	output [63:0] Sum;
	output Cout;
	input [63:0] A;
	input [63:0] B;
	input Cin;

	// define the initial block of KGP
	wire [1:0] x_00;
	assign x_00 = {2{1'b0}};

	// First let us compute the XOR-Sum of A and B
	wire [63:0] xorSum,carry;
	assign xorSum = A ^ B;

	// Define the KGP wires
	wire[1:0] x_0[63:0];
	wire[1:0] x_1[63:0];
	wire[1:0] x_2[63:0];
	wire[1:0] x_3[63:0];
	wire[1:0] x_4[63:0];
	wire[1:0] x_5[63:0];
	wire[1:0] x_6[63:0];

	// Assign the first KGP values
	assign x_0[0][0] = A[0];
	assign x_0[1][0] = A[1];
	assign x_0[2][0] = A[2];
	assign x_0[3][0] = A[3];
	assign x_0[4][0] = A[4];
	assign x_0[5][0] = A[5];
	assign x_0[6][0] = A[6];
	assign x_0[7][0] = A[7];
	assign x_0[8][0] = A[8];
	assign x_0[9][0] = A[9];
	assign x_0[10][0] = A[10];
	assign x_0[11][0] = A[11];
	assign x_0[12][0] = A[12];
	assign x_0[13][0] = A[13];
	assign x_0[14][0] = A[14];
	assign x_0[15][0] = A[15];
	assign x_0[16][0] = A[16];
	assign x_0[17][0] = A[17];
	assign x_0[18][0] = A[18];
	assign x_0[19][0] = A[19];
	assign x_0[20][0] = A[20];
	assign x_0[21][0] = A[21];
	assign x_0[22][0] = A[22];
	assign x_0[23][0] = A[23];
	assign x_0[24][0] = A[24];
	assign x_0[25][0] = A[25];
	assign x_0[26][0] = A[26];
	assign x_0[27][0] = A[27];
	assign x_0[28][0] = A[28];
	assign x_0[29][0] = A[29];
	assign x_0[30][0] = A[30];
	assign x_0[31][0] = A[31];
	assign x_0[32][0] = A[32];
	assign x_0[33][0] = A[33];
	assign x_0[34][0] = A[34];
	assign x_0[35][0] = A[35];
	assign x_0[36][0] = A[36];
	assign x_0[37][0] = A[37];
	assign x_0[38][0] = A[38];
	assign x_0[39][0] = A[39];
	assign x_0[40][0] = A[40];
	assign x_0[41][0] = A[41];
	assign x_0[42][0] = A[42];
	assign x_0[43][0] = A[43];
	assign x_0[44][0] = A[44];
	assign x_0[45][0] = A[45];
	assign x_0[46][0] = A[46];
	assign x_0[47][0] = A[47];
	assign x_0[48][0] = A[48];
	assign x_0[49][0] = A[49];
	assign x_0[50][0] = A[50];
	assign x_0[51][0] = A[51];
	assign x_0[52][0] = A[52];
	assign x_0[53][0] = A[53];
	assign x_0[54][0] = A[54];
	assign x_0[55][0] = A[55];
	assign x_0[56][0] = A[56];
	assign x_0[57][0] = A[57];
	assign x_0[58][0] = A[58];
	assign x_0[59][0] = A[59];
	assign x_0[60][0] = A[60];
	assign x_0[61][0] = A[61];
	assign x_0[62][0] = A[62];
	assign x_0[63][0] = A[63];

	assign x_0[0][1] = B[0];
	assign x_0[1][1] = B[1];
	assign x_0[2][1] = B[2];
	assign x_0[3][1] = B[3];
	assign x_0[4][1] = B[4];
	assign x_0[5][1] = B[5];
	assign x_0[6][1] = B[6];
	assign x_0[7][1] = B[7];
	assign x_0[8][1] = B[8];
	assign x_0[9][1] = B[9];
	assign x_0[10][1] = B[10];
	assign x_0[11][1] = B[11];
	assign x_0[12][1] = B[12];
	assign x_0[13][1] = B[13];
	assign x_0[14][1] = B[14];
	assign x_0[15][1] = B[15];
	assign x_0[16][1] = B[16];
	assign x_0[17][1] = B[17];
	assign x_0[18][1] = B[18];
	assign x_0[19][1] = B[19];
	assign x_0[20][1] = B[20];
	assign x_0[21][1] = B[21];
	assign x_0[22][1] = B[22];
	assign x_0[23][1] = B[23];
	assign x_0[24][1] = B[24];
	assign x_0[25][1] = B[25];
	assign x_0[26][1] = B[26];
	assign x_0[27][1] = B[27];
	assign x_0[28][1] = B[28];
	assign x_0[29][1] = B[29];
	assign x_0[30][1] = B[30];
	assign x_0[31][1] = B[31];
	assign x_0[32][1] = B[32];
	assign x_0[33][1] = B[33];
	assign x_0[34][1] = B[34];
	assign x_0[35][1] = B[35];
	assign x_0[36][1] = B[36];
	assign x_0[37][1] = B[37];
	assign x_0[38][1] = B[38];
	assign x_0[39][1] = B[39];
	assign x_0[40][1] = B[40];
	assign x_0[41][1] = B[41];
	assign x_0[42][1] = B[42];
	assign x_0[43][1] = B[43];
	assign x_0[44][1] = B[44];
	assign x_0[45][1] = B[45];
	assign x_0[46][1] = B[46];
	assign x_0[47][1] = B[47];
	assign x_0[48][1] = B[48];
	assign x_0[49][1] = B[49];
	assign x_0[50][1] = B[50];
	assign x_0[51][1] = B[51];
	assign x_0[52][1] = B[52];
	assign x_0[53][1] = B[53];
	assign x_0[54][1] = B[54];
	assign x_0[55][1] = B[55];
	assign x_0[56][1] = B[56];
	assign x_0[57][1] = B[57];
	assign x_0[58][1] = B[58];
	assign x_0[59][1] = B[59];
	assign x_0[60][1] = B[60];
	assign x_0[61][1] = B[61];
	assign x_0[62][1] = B[62];
	assign x_0[63][1] = B[63];

	// 1st Stage of KGP - Recursive Doubling
	parallelPrefixCkt p0_63(x_1[63],x_0[63],x_0[62]);
	parallelPrefixCkt p0_62(x_1[62],x_0[62],x_0[61]);
	parallelPrefixCkt p0_61(x_1[61],x_0[61],x_0[60]);
	parallelPrefixCkt p0_60(x_1[60],x_0[60],x_0[59]);
	parallelPrefixCkt p0_59(x_1[59],x_0[59],x_0[58]);
	parallelPrefixCkt p0_58(x_1[58],x_0[58],x_0[57]);
	parallelPrefixCkt p0_57(x_1[57],x_0[57],x_0[56]);
	parallelPrefixCkt p0_56(x_1[56],x_0[56],x_0[55]);
	parallelPrefixCkt p0_55(x_1[55],x_0[55],x_0[54]);
	parallelPrefixCkt p0_54(x_1[54],x_0[54],x_0[53]);
	parallelPrefixCkt p0_53(x_1[53],x_0[53],x_0[52]);
	parallelPrefixCkt p0_52(x_1[52],x_0[52],x_0[51]);
	parallelPrefixCkt p0_51(x_1[51],x_0[51],x_0[50]);
	parallelPrefixCkt p0_50(x_1[50],x_0[50],x_0[49]);
	parallelPrefixCkt p0_49(x_1[49],x_0[49],x_0[48]);
	parallelPrefixCkt p0_48(x_1[48],x_0[48],x_0[47]);
	parallelPrefixCkt p0_47(x_1[47],x_0[47],x_0[46]);
	parallelPrefixCkt p0_46(x_1[46],x_0[46],x_0[45]);
	parallelPrefixCkt p0_45(x_1[45],x_0[45],x_0[44]);
	parallelPrefixCkt p0_44(x_1[44],x_0[44],x_0[43]);
	parallelPrefixCkt p0_43(x_1[43],x_0[43],x_0[42]);
	parallelPrefixCkt p0_42(x_1[42],x_0[42],x_0[41]);
	parallelPrefixCkt p0_41(x_1[41],x_0[41],x_0[40]);
	parallelPrefixCkt p0_40(x_1[40],x_0[40],x_0[39]);
	parallelPrefixCkt p0_39(x_1[39],x_0[39],x_0[38]);
	parallelPrefixCkt p0_38(x_1[38],x_0[38],x_0[37]);
	parallelPrefixCkt p0_37(x_1[37],x_0[37],x_0[36]);
	parallelPrefixCkt p0_36(x_1[36],x_0[36],x_0[35]);
	parallelPrefixCkt p0_35(x_1[35],x_0[35],x_0[34]);
	parallelPrefixCkt p0_34(x_1[34],x_0[34],x_0[33]);
	parallelPrefixCkt p0_33(x_1[33],x_0[33],x_0[32]);
	parallelPrefixCkt p0_32(x_1[32],x_0[32],x_0[31]);
	parallelPrefixCkt p0_31(x_1[31],x_0[31],x_0[30]);
	parallelPrefixCkt p0_30(x_1[30],x_0[30],x_0[29]);
	parallelPrefixCkt p0_29(x_1[29],x_0[29],x_0[28]);
	parallelPrefixCkt p0_28(x_1[28],x_0[28],x_0[27]);
	parallelPrefixCkt p0_27(x_1[27],x_0[27],x_0[26]);
	parallelPrefixCkt p0_26(x_1[26],x_0[26],x_0[25]);
	parallelPrefixCkt p0_25(x_1[25],x_0[25],x_0[24]);
	parallelPrefixCkt p0_24(x_1[24],x_0[24],x_0[23]);
	parallelPrefixCkt p0_23(x_1[23],x_0[23],x_0[22]);
	parallelPrefixCkt p0_22(x_1[22],x_0[22],x_0[21]);
	parallelPrefixCkt p0_21(x_1[21],x_0[21],x_0[20]);
	parallelPrefixCkt p0_20(x_1[20],x_0[20],x_0[19]);
	parallelPrefixCkt p0_19(x_1[19],x_0[19],x_0[18]);
	parallelPrefixCkt p0_18(x_1[18],x_0[18],x_0[17]);
	parallelPrefixCkt p0_17(x_1[17],x_0[17],x_0[16]);
	parallelPrefixCkt p0_16(x_1[16],x_0[16],x_0[15]);
	parallelPrefixCkt p0_15(x_1[15],x_0[15],x_0[14]);
	parallelPrefixCkt p0_14(x_1[14],x_0[14],x_0[13]);
	parallelPrefixCkt p0_13(x_1[13],x_0[13],x_0[12]);
	parallelPrefixCkt p0_12(x_1[12],x_0[12],x_0[11]);
	parallelPrefixCkt p0_11(x_1[11],x_0[11],x_0[10]);
	parallelPrefixCkt p0_10(x_1[10],x_0[10],x_0[9]);
	parallelPrefixCkt p0_9(x_1[9],x_0[9],x_0[8]);
	parallelPrefixCkt p0_8(x_1[8],x_0[8],x_0[7]);
	parallelPrefixCkt p0_7(x_1[7],x_0[7],x_0[6]);
	parallelPrefixCkt p0_6(x_1[6],x_0[6],x_0[5]);
	parallelPrefixCkt p0_5(x_1[5],x_0[5],x_0[4]);
	parallelPrefixCkt p0_4(x_1[4],x_0[4],x_0[3]);
	parallelPrefixCkt p0_3(x_1[3],x_0[3],x_0[2]);
	parallelPrefixCkt p0_2(x_1[2],x_0[2],x_0[1]);
	parallelPrefixCkt p0_1(x_1[1],x_0[1],x_0[0]);
	parallelPrefixCkt p0_0(x_1[0],x_0[0],x_00);

	// 2nd stage of KGP
	parallelPrefixCkt p1_63(x_2[63],x_1[63],x_1[61]);
	parallelPrefixCkt p1_62(x_2[62],x_1[62],x_1[60]);
	parallelPrefixCkt p1_61(x_2[61],x_1[61],x_1[59]);
	parallelPrefixCkt p1_60(x_2[60],x_1[60],x_1[58]);
	parallelPrefixCkt p1_59(x_2[59],x_1[59],x_1[57]);
	parallelPrefixCkt p1_58(x_2[58],x_1[58],x_1[56]);
	parallelPrefixCkt p1_57(x_2[57],x_1[57],x_1[55]);
	parallelPrefixCkt p1_56(x_2[56],x_1[56],x_1[54]);
	parallelPrefixCkt p1_55(x_2[55],x_1[55],x_1[53]);
	parallelPrefixCkt p1_54(x_2[54],x_1[54],x_1[52]);
	parallelPrefixCkt p1_53(x_2[53],x_1[53],x_1[51]);
	parallelPrefixCkt p1_52(x_2[52],x_1[52],x_1[50]);
	parallelPrefixCkt p1_51(x_2[51],x_1[51],x_1[49]);
	parallelPrefixCkt p1_50(x_2[50],x_1[50],x_1[48]);
	parallelPrefixCkt p1_49(x_2[49],x_1[49],x_1[47]);
	parallelPrefixCkt p1_48(x_2[48],x_1[48],x_1[46]);
	parallelPrefixCkt p1_47(x_2[47],x_1[47],x_1[45]);
	parallelPrefixCkt p1_46(x_2[46],x_1[46],x_1[44]);
	parallelPrefixCkt p1_45(x_2[45],x_1[45],x_1[43]);
	parallelPrefixCkt p1_44(x_2[44],x_1[44],x_1[42]);
	parallelPrefixCkt p1_43(x_2[43],x_1[43],x_1[41]);
	parallelPrefixCkt p1_42(x_2[42],x_1[42],x_1[40]);
	parallelPrefixCkt p1_41(x_2[41],x_1[41],x_1[39]);
	parallelPrefixCkt p1_40(x_2[40],x_1[40],x_1[38]);
	parallelPrefixCkt p1_39(x_2[39],x_1[39],x_1[37]);
	parallelPrefixCkt p1_38(x_2[38],x_1[38],x_1[36]);
	parallelPrefixCkt p1_37(x_2[37],x_1[37],x_1[35]);
	parallelPrefixCkt p1_36(x_2[36],x_1[36],x_1[34]);
	parallelPrefixCkt p1_35(x_2[35],x_1[35],x_1[33]);
	parallelPrefixCkt p1_34(x_2[34],x_1[34],x_1[32]);
	parallelPrefixCkt p1_33(x_2[33],x_1[33],x_1[31]);
	parallelPrefixCkt p1_32(x_2[32],x_1[32],x_1[30]);
	parallelPrefixCkt p1_31(x_2[31],x_1[31],x_1[29]);
	parallelPrefixCkt p1_30(x_2[30],x_1[30],x_1[28]);
	parallelPrefixCkt p1_29(x_2[29],x_1[29],x_1[27]);
	parallelPrefixCkt p1_28(x_2[28],x_1[28],x_1[26]);
	parallelPrefixCkt p1_27(x_2[27],x_1[27],x_1[25]);
	parallelPrefixCkt p1_26(x_2[26],x_1[26],x_1[24]);
	parallelPrefixCkt p1_25(x_2[25],x_1[25],x_1[23]);
	parallelPrefixCkt p1_24(x_2[24],x_1[24],x_1[22]);
	parallelPrefixCkt p1_23(x_2[23],x_1[23],x_1[21]);
	parallelPrefixCkt p1_22(x_2[22],x_1[22],x_1[20]);
	parallelPrefixCkt p1_21(x_2[21],x_1[21],x_1[19]);
	parallelPrefixCkt p1_20(x_2[20],x_1[20],x_1[18]);
	parallelPrefixCkt p1_19(x_2[19],x_1[19],x_1[17]);
	parallelPrefixCkt p1_18(x_2[18],x_1[18],x_1[16]);
	parallelPrefixCkt p1_17(x_2[17],x_1[17],x_1[15]);
	parallelPrefixCkt p1_16(x_2[16],x_1[16],x_1[14]);
	parallelPrefixCkt p1_15(x_2[15],x_1[15],x_1[13]);
	parallelPrefixCkt p1_14(x_2[14],x_1[14],x_1[12]);
	parallelPrefixCkt p1_13(x_2[13],x_1[13],x_1[11]);
	parallelPrefixCkt p1_12(x_2[12],x_1[12],x_1[10]);
	parallelPrefixCkt p1_11(x_2[11],x_1[11],x_1[9]);
	parallelPrefixCkt p1_10(x_2[10],x_1[10],x_1[8]);
	parallelPrefixCkt p1_9(x_2[9],x_1[9],x_1[7]);
	parallelPrefixCkt p1_8(x_2[8],x_1[8],x_1[6]);
	parallelPrefixCkt p1_7(x_2[7],x_1[7],x_1[5]);
	parallelPrefixCkt p1_6(x_2[6],x_1[6],x_1[4]);
	parallelPrefixCkt p1_5(x_2[5],x_1[5],x_1[3]);
	parallelPrefixCkt p1_4(x_2[4],x_1[4],x_1[2]);
	parallelPrefixCkt p1_3(x_2[3],x_1[3],x_1[1]);
	parallelPrefixCkt p1_2(x_2[2],x_1[2],x_1[0]);
	parallelPrefixCkt p1_1(x_2[1],x_1[1],x_00);
	parallelPrefixCkt p1_0(x_2[0],x_1[0],x_00);

	// 3rd stage of KGP
	parallelPrefixCkt p2_63(x_3[63],x_2[63],x_2[59]);
	parallelPrefixCkt p2_62(x_3[62],x_2[62],x_2[58]);
	parallelPrefixCkt p2_61(x_3[61],x_2[61],x_2[57]);
	parallelPrefixCkt p2_60(x_3[60],x_2[60],x_2[56]);
	parallelPrefixCkt p2_59(x_3[59],x_2[59],x_2[55]);
	parallelPrefixCkt p2_58(x_3[58],x_2[58],x_2[54]);
	parallelPrefixCkt p2_57(x_3[57],x_2[57],x_2[53]);
	parallelPrefixCkt p2_56(x_3[56],x_2[56],x_2[52]);
	parallelPrefixCkt p2_55(x_3[55],x_2[55],x_2[51]);
	parallelPrefixCkt p2_54(x_3[54],x_2[54],x_2[50]);
	parallelPrefixCkt p2_53(x_3[53],x_2[53],x_2[49]);
	parallelPrefixCkt p2_52(x_3[52],x_2[52],x_2[48]);
	parallelPrefixCkt p2_51(x_3[51],x_2[51],x_2[47]);
	parallelPrefixCkt p2_50(x_3[50],x_2[50],x_2[46]);
	parallelPrefixCkt p2_49(x_3[49],x_2[49],x_2[45]);
	parallelPrefixCkt p2_48(x_3[48],x_2[48],x_2[44]);
	parallelPrefixCkt p2_47(x_3[47],x_2[47],x_2[43]);
	parallelPrefixCkt p2_46(x_3[46],x_2[46],x_2[42]);
	parallelPrefixCkt p2_45(x_3[45],x_2[45],x_2[41]);
	parallelPrefixCkt p2_44(x_3[44],x_2[44],x_2[40]);
	parallelPrefixCkt p2_43(x_3[43],x_2[43],x_2[39]);
	parallelPrefixCkt p2_42(x_3[42],x_2[42],x_2[38]);
	parallelPrefixCkt p2_41(x_3[41],x_2[41],x_2[37]);
	parallelPrefixCkt p2_40(x_3[40],x_2[40],x_2[36]);
	parallelPrefixCkt p2_39(x_3[39],x_2[39],x_2[35]);
	parallelPrefixCkt p2_38(x_3[38],x_2[38],x_2[34]);
	parallelPrefixCkt p2_37(x_3[37],x_2[37],x_2[33]);
	parallelPrefixCkt p2_36(x_3[36],x_2[36],x_2[32]);
	parallelPrefixCkt p2_35(x_3[35],x_2[35],x_2[31]);
	parallelPrefixCkt p2_34(x_3[34],x_2[34],x_2[30]);
	parallelPrefixCkt p2_33(x_3[33],x_2[33],x_2[29]);
	parallelPrefixCkt p2_32(x_3[32],x_2[32],x_2[28]);
	parallelPrefixCkt p2_31(x_3[31],x_2[31],x_2[27]);
	parallelPrefixCkt p2_30(x_3[30],x_2[30],x_2[26]);
	parallelPrefixCkt p2_29(x_3[29],x_2[29],x_2[25]);
	parallelPrefixCkt p2_28(x_3[28],x_2[28],x_2[24]);
	parallelPrefixCkt p2_27(x_3[27],x_2[27],x_2[23]);
	parallelPrefixCkt p2_26(x_3[26],x_2[26],x_2[22]);
	parallelPrefixCkt p2_25(x_3[25],x_2[25],x_2[21]);
	parallelPrefixCkt p2_24(x_3[24],x_2[24],x_2[20]);
	parallelPrefixCkt p2_23(x_3[23],x_2[23],x_2[19]);
	parallelPrefixCkt p2_22(x_3[22],x_2[22],x_2[18]);
	parallelPrefixCkt p2_21(x_3[21],x_2[21],x_2[17]);
	parallelPrefixCkt p2_20(x_3[20],x_2[20],x_2[16]);
	parallelPrefixCkt p2_19(x_3[19],x_2[19],x_2[15]);
	parallelPrefixCkt p2_18(x_3[18],x_2[18],x_2[14]);
	parallelPrefixCkt p2_17(x_3[17],x_2[17],x_2[13]);
	parallelPrefixCkt p2_16(x_3[16],x_2[16],x_2[12]);
	parallelPrefixCkt p2_15(x_3[15],x_2[15],x_2[11]);
	parallelPrefixCkt p2_14(x_3[14],x_2[14],x_2[10]);
	parallelPrefixCkt p2_13(x_3[13],x_2[13],x_2[9]);
	parallelPrefixCkt p2_12(x_3[12],x_2[12],x_2[8]);
	parallelPrefixCkt p2_11(x_3[11],x_2[11],x_2[7]);
	parallelPrefixCkt p2_10(x_3[10],x_2[10],x_2[6]);
	parallelPrefixCkt p2_9(x_3[9],x_2[9],x_2[5]);
	parallelPrefixCkt p2_8(x_3[8],x_2[8],x_2[4]);
	parallelPrefixCkt p2_7(x_3[7],x_2[7],x_2[3]);
	parallelPrefixCkt p2_6(x_3[6],x_2[6],x_2[2]);
	parallelPrefixCkt p2_5(x_3[5],x_2[5],x_2[1]);
	parallelPrefixCkt p2_4(x_3[4],x_2[4],x_2[0]);
	parallelPrefixCkt p2_3(x_3[3],x_2[3],x_00);
	parallelPrefixCkt p2_2(x_3[2],x_2[2],x_00);
	parallelPrefixCkt p2_1(x_3[1],x_2[1],x_00);
	parallelPrefixCkt p2_0(x_3[0],x_2[0],x_00);

	// 4th stage of KGP
	parallelPrefixCkt p3_63(x_4[63],x_3[63],x_3[55]);
	parallelPrefixCkt p3_62(x_4[62],x_3[62],x_3[54]);
	parallelPrefixCkt p3_61(x_4[61],x_3[61],x_3[53]);
	parallelPrefixCkt p3_60(x_4[60],x_3[60],x_3[52]);
	parallelPrefixCkt p3_59(x_4[59],x_3[59],x_3[51]);
	parallelPrefixCkt p3_58(x_4[58],x_3[58],x_3[50]);
	parallelPrefixCkt p3_57(x_4[57],x_3[57],x_3[49]);
	parallelPrefixCkt p3_56(x_4[56],x_3[56],x_3[48]);
	parallelPrefixCkt p3_55(x_4[55],x_3[55],x_3[47]);
	parallelPrefixCkt p3_54(x_4[54],x_3[54],x_3[46]);
	parallelPrefixCkt p3_53(x_4[53],x_3[53],x_3[45]);
	parallelPrefixCkt p3_52(x_4[52],x_3[52],x_3[44]);
	parallelPrefixCkt p3_51(x_4[51],x_3[51],x_3[43]);
	parallelPrefixCkt p3_50(x_4[50],x_3[50],x_3[42]);
	parallelPrefixCkt p3_49(x_4[49],x_3[49],x_3[41]);
	parallelPrefixCkt p3_48(x_4[48],x_3[48],x_3[40]);
	parallelPrefixCkt p3_47(x_4[47],x_3[47],x_3[39]);
	parallelPrefixCkt p3_46(x_4[46],x_3[46],x_3[38]);
	parallelPrefixCkt p3_45(x_4[45],x_3[45],x_3[37]);
	parallelPrefixCkt p3_44(x_4[44],x_3[44],x_3[36]);
	parallelPrefixCkt p3_43(x_4[43],x_3[43],x_3[35]);
	parallelPrefixCkt p3_42(x_4[42],x_3[42],x_3[34]);
	parallelPrefixCkt p3_41(x_4[41],x_3[41],x_3[33]);
	parallelPrefixCkt p3_40(x_4[40],x_3[40],x_3[32]);
	parallelPrefixCkt p3_39(x_4[39],x_3[39],x_3[31]);
	parallelPrefixCkt p3_38(x_4[38],x_3[38],x_3[30]);
	parallelPrefixCkt p3_37(x_4[37],x_3[37],x_3[29]);
	parallelPrefixCkt p3_36(x_4[36],x_3[36],x_3[28]);
	parallelPrefixCkt p3_35(x_4[35],x_3[35],x_3[27]);
	parallelPrefixCkt p3_34(x_4[34],x_3[34],x_3[26]);
	parallelPrefixCkt p3_33(x_4[33],x_3[33],x_3[25]);
	parallelPrefixCkt p3_32(x_4[32],x_3[32],x_3[24]);
	parallelPrefixCkt p3_31(x_4[31],x_3[31],x_3[23]);
	parallelPrefixCkt p3_30(x_4[30],x_3[30],x_3[22]);
	parallelPrefixCkt p3_29(x_4[29],x_3[29],x_3[21]);
	parallelPrefixCkt p3_28(x_4[28],x_3[28],x_3[20]);
	parallelPrefixCkt p3_27(x_4[27],x_3[27],x_3[19]);
	parallelPrefixCkt p3_26(x_4[26],x_3[26],x_3[18]);
	parallelPrefixCkt p3_25(x_4[25],x_3[25],x_3[17]);
	parallelPrefixCkt p3_24(x_4[24],x_3[24],x_3[16]);
	parallelPrefixCkt p3_23(x_4[23],x_3[23],x_3[15]);
	parallelPrefixCkt p3_22(x_4[22],x_3[22],x_3[14]);
	parallelPrefixCkt p3_21(x_4[21],x_3[21],x_3[13]);
	parallelPrefixCkt p3_20(x_4[20],x_3[20],x_3[12]);
	parallelPrefixCkt p3_19(x_4[19],x_3[19],x_3[11]);
	parallelPrefixCkt p3_18(x_4[18],x_3[18],x_3[10]);
	parallelPrefixCkt p3_17(x_4[17],x_3[17],x_3[9]);
	parallelPrefixCkt p3_16(x_4[16],x_3[16],x_3[8]);
	parallelPrefixCkt p3_15(x_4[15],x_3[15],x_3[7]);
	parallelPrefixCkt p3_14(x_4[14],x_3[14],x_3[6]);
	parallelPrefixCkt p3_13(x_4[13],x_3[13],x_3[5]);
	parallelPrefixCkt p3_12(x_4[12],x_3[12],x_3[4]);
	parallelPrefixCkt p3_11(x_4[11],x_3[11],x_3[3]);
	parallelPrefixCkt p3_10(x_4[10],x_3[10],x_3[2]);
	parallelPrefixCkt p3_9(x_4[9],x_3[9],x_3[1]);
	parallelPrefixCkt p3_8(x_4[8],x_3[8],x_3[0]);
	parallelPrefixCkt p3_7(x_4[7],x_3[7],x_00);
	parallelPrefixCkt p3_6(x_4[6],x_3[6],x_00);
	parallelPrefixCkt p3_5(x_4[5],x_3[5],x_00);
	parallelPrefixCkt p3_4(x_4[4],x_3[4],x_00);
	parallelPrefixCkt p3_3(x_4[3],x_3[3],x_00);
	parallelPrefixCkt p3_2(x_4[2],x_3[2],x_00);
	parallelPrefixCkt p3_1(x_4[1],x_3[1],x_00);
	parallelPrefixCkt p3_0(x_4[0],x_3[0],x_00);

	// 5th stage of KGP
	parallelPrefixCkt p4_63(x_5[63],x_4[63],x_4[47]);
	parallelPrefixCkt p4_62(x_5[62],x_4[62],x_4[46]);
	parallelPrefixCkt p4_61(x_5[61],x_4[61],x_4[45]);
	parallelPrefixCkt p4_60(x_5[60],x_4[60],x_4[44]);
	parallelPrefixCkt p4_59(x_5[59],x_4[59],x_4[43]);
	parallelPrefixCkt p4_58(x_5[58],x_4[58],x_4[42]);
	parallelPrefixCkt p4_57(x_5[57],x_4[57],x_4[41]);
	parallelPrefixCkt p4_56(x_5[56],x_4[56],x_4[40]);
	parallelPrefixCkt p4_55(x_5[55],x_4[55],x_4[39]);
	parallelPrefixCkt p4_54(x_5[54],x_4[54],x_4[38]);
	parallelPrefixCkt p4_53(x_5[53],x_4[53],x_4[37]);
	parallelPrefixCkt p4_52(x_5[52],x_4[52],x_4[36]);
	parallelPrefixCkt p4_51(x_5[51],x_4[51],x_4[35]);
	parallelPrefixCkt p4_50(x_5[50],x_4[50],x_4[34]);
	parallelPrefixCkt p4_49(x_5[49],x_4[49],x_4[33]);
	parallelPrefixCkt p4_48(x_5[48],x_4[48],x_4[32]);
	parallelPrefixCkt p4_47(x_5[47],x_4[47],x_4[31]);
	parallelPrefixCkt p4_46(x_5[46],x_4[46],x_4[30]);
	parallelPrefixCkt p4_45(x_5[45],x_4[45],x_4[29]);
	parallelPrefixCkt p4_44(x_5[44],x_4[44],x_4[28]);
	parallelPrefixCkt p4_43(x_5[43],x_4[43],x_4[27]);
	parallelPrefixCkt p4_42(x_5[42],x_4[42],x_4[26]);
	parallelPrefixCkt p4_41(x_5[41],x_4[41],x_4[25]);
	parallelPrefixCkt p4_40(x_5[40],x_4[40],x_4[24]);
	parallelPrefixCkt p4_39(x_5[39],x_4[39],x_4[23]);
	parallelPrefixCkt p4_38(x_5[38],x_4[38],x_4[22]);
	parallelPrefixCkt p4_37(x_5[37],x_4[37],x_4[21]);
	parallelPrefixCkt p4_36(x_5[36],x_4[36],x_4[20]);
	parallelPrefixCkt p4_35(x_5[35],x_4[35],x_4[19]);
	parallelPrefixCkt p4_34(x_5[34],x_4[34],x_4[18]);
	parallelPrefixCkt p4_33(x_5[33],x_4[33],x_4[17]);
	parallelPrefixCkt p4_32(x_5[32],x_4[32],x_4[16]);
	parallelPrefixCkt p4_31(x_5[31],x_4[31],x_4[15]);
	parallelPrefixCkt p4_30(x_5[30],x_4[30],x_4[14]);
	parallelPrefixCkt p4_29(x_5[29],x_4[29],x_4[13]);
	parallelPrefixCkt p4_28(x_5[28],x_4[28],x_4[12]);
	parallelPrefixCkt p4_27(x_5[27],x_4[27],x_4[11]);
	parallelPrefixCkt p4_26(x_5[26],x_4[26],x_4[10]);
	parallelPrefixCkt p4_25(x_5[25],x_4[25],x_4[9]);
	parallelPrefixCkt p4_24(x_5[24],x_4[24],x_4[8]);
	parallelPrefixCkt p4_23(x_5[23],x_4[23],x_4[7]);
	parallelPrefixCkt p4_22(x_5[22],x_4[22],x_4[6]);
	parallelPrefixCkt p4_21(x_5[21],x_4[21],x_4[5]);
	parallelPrefixCkt p4_20(x_5[20],x_4[20],x_4[4]);
	parallelPrefixCkt p4_19(x_5[19],x_4[19],x_4[3]);
	parallelPrefixCkt p4_18(x_5[18],x_4[18],x_4[2]);
	parallelPrefixCkt p4_17(x_5[17],x_4[17],x_4[1]);
	parallelPrefixCkt p4_16(x_5[16],x_4[16],x_4[0]);
	parallelPrefixCkt p4_15(x_5[15],x_4[15],x_00);
	parallelPrefixCkt p4_14(x_5[14],x_4[14],x_00);
	parallelPrefixCkt p4_13(x_5[13],x_4[13],x_00);
	parallelPrefixCkt p4_12(x_5[12],x_4[12],x_00);
	parallelPrefixCkt p4_11(x_5[11],x_4[11],x_00);
	parallelPrefixCkt p4_10(x_5[10],x_4[10],x_00);
	parallelPrefixCkt p4_9(x_5[9],x_4[9],x_00);
	parallelPrefixCkt p4_8(x_5[8],x_4[8],x_00);
	parallelPrefixCkt p4_7(x_5[7],x_4[7],x_00);
	parallelPrefixCkt p4_6(x_5[6],x_4[6],x_00);
	parallelPrefixCkt p4_5(x_5[5],x_4[5],x_00);
	parallelPrefixCkt p4_4(x_5[4],x_4[4],x_00);
	parallelPrefixCkt p4_3(x_5[3],x_4[3],x_00);
	parallelPrefixCkt p4_2(x_5[2],x_4[2],x_00);
	parallelPrefixCkt p4_1(x_5[1],x_4[1],x_00);
	parallelPrefixCkt p4_0(x_5[0],x_4[0],x_00);

	// 6th stage
	parallelPrefixCkt p5_63(x_6[63],x_5[63],x_5[31]);
	parallelPrefixCkt p5_62(x_6[62],x_5[62],x_5[30]);
	parallelPrefixCkt p5_61(x_6[61],x_5[61],x_5[29]);
	parallelPrefixCkt p5_60(x_6[60],x_5[60],x_5[28]);
	parallelPrefixCkt p5_59(x_6[59],x_5[59],x_5[27]);
	parallelPrefixCkt p5_58(x_6[58],x_5[58],x_5[26]);
	parallelPrefixCkt p5_57(x_6[57],x_5[57],x_5[25]);
	parallelPrefixCkt p5_56(x_6[56],x_5[56],x_5[24]);
	parallelPrefixCkt p5_55(x_6[55],x_5[55],x_5[23]);
	parallelPrefixCkt p5_54(x_6[54],x_5[54],x_5[22]);
	parallelPrefixCkt p5_53(x_6[53],x_5[53],x_5[21]);
	parallelPrefixCkt p5_52(x_6[52],x_5[52],x_5[20]);
	parallelPrefixCkt p5_51(x_6[51],x_5[51],x_5[19]);
	parallelPrefixCkt p5_50(x_6[50],x_5[50],x_5[18]);
	parallelPrefixCkt p5_49(x_6[49],x_5[49],x_5[17]);
	parallelPrefixCkt p5_48(x_6[48],x_5[48],x_5[16]);
	parallelPrefixCkt p5_47(x_6[47],x_5[47],x_5[15]);
	parallelPrefixCkt p5_46(x_6[46],x_5[46],x_5[14]);
	parallelPrefixCkt p5_45(x_6[45],x_5[45],x_5[13]);
	parallelPrefixCkt p5_44(x_6[44],x_5[44],x_5[12]);
	parallelPrefixCkt p5_43(x_6[43],x_5[43],x_5[11]);
	parallelPrefixCkt p5_42(x_6[42],x_5[42],x_5[10]);
	parallelPrefixCkt p5_41(x_6[41],x_5[41],x_5[9]);
	parallelPrefixCkt p5_40(x_6[40],x_5[40],x_5[8]);
	parallelPrefixCkt p5_39(x_6[39],x_5[39],x_5[7]);
	parallelPrefixCkt p5_38(x_6[38],x_5[38],x_5[6]);
	parallelPrefixCkt p5_37(x_6[37],x_5[37],x_5[5]);
	parallelPrefixCkt p5_36(x_6[36],x_5[36],x_5[4]);
	parallelPrefixCkt p5_35(x_6[35],x_5[35],x_5[3]);
	parallelPrefixCkt p5_34(x_6[34],x_5[34],x_5[2]);
	parallelPrefixCkt p5_33(x_6[33],x_5[33],x_5[1]);
	parallelPrefixCkt p5_32(x_6[32],x_5[32],x_5[0]);
	parallelPrefixCkt p5_31(x_6[31],x_5[31],x_00);
	parallelPrefixCkt p5_30(x_6[30],x_5[30],x_00);
	parallelPrefixCkt p5_29(x_6[29],x_5[29],x_00);
	parallelPrefixCkt p5_28(x_6[28],x_5[28],x_00);
	parallelPrefixCkt p5_27(x_6[27],x_5[27],x_00);
	parallelPrefixCkt p5_26(x_6[26],x_5[26],x_00);
	parallelPrefixCkt p5_25(x_6[25],x_5[25],x_00);
	parallelPrefixCkt p5_24(x_6[24],x_5[24],x_00);
	parallelPrefixCkt p5_23(x_6[23],x_5[23],x_00);
	parallelPrefixCkt p5_22(x_6[22],x_5[22],x_00);
	parallelPrefixCkt p5_21(x_6[21],x_5[21],x_00);
	parallelPrefixCkt p5_20(x_6[20],x_5[20],x_00);
	parallelPrefixCkt p5_19(x_6[19],x_5[19],x_00);
	parallelPrefixCkt p5_18(x_6[18],x_5[18],x_00);
	parallelPrefixCkt p5_17(x_6[17],x_5[17],x_00);
	parallelPrefixCkt p5_16(x_6[16],x_5[16],x_00);
	parallelPrefixCkt p5_15(x_6[15],x_5[15],x_00);
	parallelPrefixCkt p5_14(x_6[14],x_5[14],x_00);
	parallelPrefixCkt p5_13(x_6[13],x_5[13],x_00);
	parallelPrefixCkt p5_12(x_6[12],x_5[12],x_00);
	parallelPrefixCkt p5_11(x_6[11],x_5[11],x_00);
	parallelPrefixCkt p5_10(x_6[10],x_5[10],x_00);
	parallelPrefixCkt p5_9(x_6[9],x_5[9],x_00);
	parallelPrefixCkt p5_8(x_6[8],x_5[8],x_00);
	parallelPrefixCkt p5_7(x_6[7],x_5[7],x_00);
	parallelPrefixCkt p5_6(x_6[6],x_5[6],x_00);
	parallelPrefixCkt p5_5(x_6[5],x_5[5],x_00);
	parallelPrefixCkt p5_4(x_6[4],x_5[4],x_00);
	parallelPrefixCkt p5_3(x_6[3],x_5[3],x_00);
	parallelPrefixCkt p5_2(x_6[2],x_5[2],x_00);
	parallelPrefixCkt p5_1(x_6[1],x_5[1],x_00);
	parallelPrefixCkt p5_0(x_6[0],x_5[0],x_00);



	// MSB of last stage KGP is carry
	assign carry[0] = x_6[0][0];
	assign carry[1] = x_6[1][0];
	assign carry[2] = x_6[2][0];
	assign carry[3] = x_6[3][0];
	assign carry[4] = x_6[4][0];
	assign carry[5] = x_6[5][0];
	assign carry[6] = x_6[6][0];
	assign carry[7] = x_6[7][0];
	assign carry[8] = x_6[8][0];
	assign carry[9] = x_6[9][0];
	assign carry[10] = x_6[10][0];
	assign carry[11] = x_6[11][0];
	assign carry[12] = x_6[12][0];
	assign carry[13] = x_6[13][0];
	assign carry[14] = x_6[14][0];
	assign carry[15] = x_6[15][0];
	assign carry[16] = x_6[16][0];
	assign carry[17] = x_6[17][0];
	assign carry[18] = x_6[18][0];
	assign carry[19] = x_6[19][0];
	assign carry[20] = x_6[20][0];
	assign carry[21] = x_6[21][0];
	assign carry[22] = x_6[22][0];
	assign carry[23] = x_6[23][0];
	assign carry[24] = x_6[24][0];
	assign carry[25] = x_6[25][0];
	assign carry[26] = x_6[26][0];
	assign carry[27] = x_6[27][0];
	assign carry[28] = x_6[28][0];
	assign carry[29] = x_6[29][0];
	assign carry[30] = x_6[30][0];
	assign carry[31] = x_6[31][0];
	assign carry[32] = x_6[32][0];
	assign carry[33] = x_6[33][0];
	assign carry[34] = x_6[34][0];
	assign carry[35] = x_6[35][0];
	assign carry[36] = x_6[36][0];
	assign carry[37] = x_6[37][0];
	assign carry[38] = x_6[38][0];
	assign carry[39] = x_6[39][0];
	assign carry[40] = x_6[40][0];
	assign carry[41] = x_6[41][0];
	assign carry[42] = x_6[42][0];
	assign carry[43] = x_6[43][0];
	assign carry[44] = x_6[44][0];
	assign carry[45] = x_6[45][0];
	assign carry[46] = x_6[46][0];
	assign carry[47] = x_6[47][0];
	assign carry[48] = x_6[48][0];
	assign carry[49] = x_6[49][0];
	assign carry[50] = x_6[50][0];
	assign carry[51] = x_6[51][0];
	assign carry[52] = x_6[52][0];
	assign carry[53] = x_6[53][0];
	assign carry[54] = x_6[54][0];
	assign carry[55] = x_6[55][0];
	assign carry[56] = x_6[56][0];
	assign carry[57] = x_6[57][0];
	assign carry[58] = x_6[58][0];
	assign carry[59] = x_6[59][0];
	assign carry[60] = x_6[60][0];
	assign carry[61] = x_6[61][0];
	assign carry[62] = x_6[62][0];
	assign carry[63] = x_6[63][0];

	// Compute Sum
	assign Sum[0] = xorSum[0];
	assign Sum[1] = xorSum[1] ^ carry[0];
	assign Sum[2] = xorSum[2] ^ carry[1];
	assign Sum[3] = xorSum[3] ^ carry[2];
	assign Sum[4] = xorSum[4] ^ carry[3];
	assign Sum[5] = xorSum[5] ^ carry[4];
	assign Sum[6] = xorSum[6] ^ carry[5];
	assign Sum[7] = xorSum[7] ^ carry[6];
	assign Sum[8] = xorSum[8] ^ carry[7];
	assign Sum[9] = xorSum[9] ^ carry[8];
	assign Sum[10] = xorSum[10] ^ carry[9];
	assign Sum[11] = xorSum[11] ^ carry[10];
	assign Sum[12] = xorSum[12] ^ carry[11];
	assign Sum[13] = xorSum[13] ^ carry[12];
	assign Sum[14] = xorSum[14] ^ carry[13];
	assign Sum[15] = xorSum[15] ^ carry[14];
	assign Sum[16] = xorSum[16] ^ carry[15];
	assign Sum[17] = xorSum[17] ^ carry[16];
	assign Sum[18] = xorSum[18] ^ carry[17];
	assign Sum[19] = xorSum[19] ^ carry[18];
	assign Sum[20] = xorSum[20] ^ carry[19];
	assign Sum[21] = xorSum[21] ^ carry[20];
	assign Sum[22] = xorSum[22] ^ carry[21];
	assign Sum[23] = xorSum[23] ^ carry[22];
	assign Sum[24] = xorSum[24] ^ carry[23];
	assign Sum[25] = xorSum[25] ^ carry[24];
	assign Sum[26] = xorSum[26] ^ carry[25];
	assign Sum[27] = xorSum[27] ^ carry[26];
	assign Sum[28] = xorSum[28] ^ carry[27];
	assign Sum[29] = xorSum[29] ^ carry[28];
	assign Sum[30] = xorSum[30] ^ carry[29];
	assign Sum[31] = xorSum[31] ^ carry[30];
	assign Sum[32] = xorSum[32] ^ carry[31];
	assign Sum[33] = xorSum[33] ^ carry[32];
	assign Sum[34] = xorSum[34] ^ carry[33];
	assign Sum[35] = xorSum[35] ^ carry[34];
	assign Sum[36] = xorSum[36] ^ carry[35];
	assign Sum[37] = xorSum[37] ^ carry[36];
	assign Sum[38] = xorSum[38] ^ carry[37];
	assign Sum[39] = xorSum[39] ^ carry[38];
	assign Sum[40] = xorSum[40] ^ carry[39];
	assign Sum[41] = xorSum[41] ^ carry[40];
	assign Sum[42] = xorSum[42] ^ carry[41];
	assign Sum[43] = xorSum[43] ^ carry[42];
	assign Sum[44] = xorSum[44] ^ carry[43];
	assign Sum[45] = xorSum[45] ^ carry[44];
	assign Sum[46] = xorSum[46] ^ carry[45];
	assign Sum[47] = xorSum[47] ^ carry[46];
	assign Sum[48] = xorSum[48] ^ carry[47];
	assign Sum[49] = xorSum[49] ^ carry[48];
	assign Sum[50] = xorSum[50] ^ carry[49];
	assign Sum[51] = xorSum[51] ^ carry[50];
	assign Sum[52] = xorSum[52] ^ carry[51];
	assign Sum[53] = xorSum[53] ^ carry[52];
	assign Sum[54] = xorSum[54] ^ carry[53];
	assign Sum[55] = xorSum[55] ^ carry[54];
	assign Sum[56] = xorSum[56] ^ carry[55];
	assign Sum[57] = xorSum[57] ^ carry[56];
	assign Sum[58] = xorSum[58] ^ carry[57];
	assign Sum[59] = xorSum[59] ^ carry[58];
	assign Sum[60] = xorSum[60] ^ carry[59];
	assign Sum[61] = xorSum[61] ^ carry[60];
	assign Sum[62] = xorSum[62] ^ carry[61];
	assign Sum[63] = xorSum[63] ^ carry[62];
    assign Cout = carry[63];

endmodule