`include "fpAdd.v"

module top;
	reg[31:0] X1,X2;
	wire[31:0] X3;

	fpADD_32 fp_0 (X3 ,X1, X2);

	// Setup the monitoring for the signal values
	initial
	begin
		$monitor($time," X1 = %b,  X2 = %b --- X3 = %b\n",X1,X2,X3);
		$dumpfile("fpa.vcd");
		$dumpvars;
	end

	// Simulate the inputs
	initial
	begin
		X1 = 0; X2 = 0;

		#5 X2 = 32'b01000001000111000000000000000000; X1 = 32'b00111111000100000000000000000000;

		#5 X2 = 32'b01000000100000000000000000000000; X1 = 32'b00111101110011001100110011001101;

		#5 X1 = 32'b01000000100000000000000000000000; X2 = 32'b10111110100000000000000000000000;

		#5 X1 = 32'b01000000100001000010100011110110; X2 = 32'b01000000000110011001100110011010;

		#5 X1 = 32'b11000000100000000000000000000000; X2 = 32'b00111110100000000000000000000000;

		#5 X1 = 32'b01000000100000000000000000000000; X2 = 32'b11000000110010000000000000000000;

		#5 X1 = 32'b01000000100000000000000000000000; X2 = 32'b11000000100000000000000000000000;

		// -4 + (-4.0078125)
		#5 X1 = 32'b11000000100000000000000000000000; X2 = 32'b11000000100000000100000000000000;

		// -2312.12 + (-142.912)
		#5 X1 = 32'b11000101000100001000000111101100; X2 = 32'b11000011000011101110100101111001;
		
		// -990.99 + 0.99
		#5 X1 = 32'b11000100011101111011111101011100; X2 = 32'b00111111011111010111000010100100;

		//  inf  + 3
		#5 X1 = 32'b01111111100000000000000000000000; X2 = 32'b01000000010000000000000000000000;
	end

endmodule