`include "multiplexers.v"

module logicUnit(Y, X1, X2, opcode);

	// I/O Port Declarations
	output[31:0] Y;
	input[31:0] X1,X2;
	input[2:0] opcode;

	// Get the result of the 8 logical operations onto an 8 32 bit wide wire
	wire[31:0] Z[7:0];
	assign Z[0] = X1 & X2;
	assign Z[1] = X1 ^ X2;
	assign Z[2] = X1 ~& X2;
	assign Z[3] = X1 | X2;
	assign Z[4] = ~X1;
	assign Z[5] = X1 ~| X2;
	assign Z[6] = ~X1 + 1'b1;
	assign Z[7] = X1 ~^ X2;
	
	// Define 32 8:1 MUXES to get the output
	mux_8_1 m_0(Y[0],{Z[7][0],Z[6][0],Z[5][0],Z[4][0],Z[3][0],Z[2][0],Z[1][0],Z[0][0]},opcode);
	mux_8_1 m_1(Y[1],{Z[7][1],Z[6][1],Z[5][1],Z[4][1],Z[3][1],Z[2][1],Z[1][1],Z[0][1]},opcode);
	mux_8_1 m_2(Y[2],{Z[7][2],Z[6][2],Z[5][2],Z[4][2],Z[3][2],Z[2][2],Z[1][2],Z[0][2]},opcode);
	mux_8_1 m_3(Y[3],{Z[7][3],Z[6][3],Z[5][3],Z[4][3],Z[3][3],Z[2][3],Z[1][3],Z[0][3]},opcode);
	mux_8_1 m_4(Y[4],{Z[7][4],Z[6][4],Z[5][4],Z[4][4],Z[3][4],Z[2][4],Z[1][4],Z[0][4]},opcode);
	mux_8_1 m_5(Y[5],{Z[7][5],Z[6][5],Z[5][5],Z[4][5],Z[3][5],Z[2][5],Z[1][5],Z[0][5]},opcode);
	mux_8_1 m_6(Y[6],{Z[7][6],Z[6][6],Z[5][6],Z[4][6],Z[3][6],Z[2][6],Z[1][6],Z[0][6]},opcode);
	mux_8_1 m_7(Y[7],{Z[7][7],Z[6][7],Z[5][7],Z[4][7],Z[3][7],Z[2][7],Z[1][7],Z[0][7]},opcode);
	mux_8_1 m_8(Y[8],{Z[7][8],Z[6][8],Z[5][8],Z[4][8],Z[3][8],Z[2][8],Z[1][8],Z[0][8]},opcode);
	mux_8_1 m_9(Y[9],{Z[7][9],Z[6][9],Z[5][9],Z[4][9],Z[3][9],Z[2][9],Z[1][9],Z[0][9]},opcode);
	mux_8_1 m_10(Y[10],{Z[7][10],Z[6][10],Z[5][10],Z[4][10],Z[3][10],Z[2][10],Z[1][10],Z[0][10]},opcode);
	mux_8_1 m_11(Y[11],{Z[7][11],Z[6][11],Z[5][11],Z[4][11],Z[3][11],Z[2][11],Z[1][11],Z[0][11]},opcode);
	mux_8_1 m_12(Y[12],{Z[7][12],Z[6][12],Z[5][12],Z[4][12],Z[3][12],Z[2][12],Z[1][12],Z[0][12]},opcode);
	mux_8_1 m_13(Y[13],{Z[7][13],Z[6][13],Z[5][13],Z[4][13],Z[3][13],Z[2][13],Z[1][13],Z[0][13]},opcode);
	mux_8_1 m_14(Y[14],{Z[7][14],Z[6][14],Z[5][14],Z[4][14],Z[3][14],Z[2][14],Z[1][14],Z[0][14]},opcode);
	mux_8_1 m_15(Y[15],{Z[7][15],Z[6][15],Z[5][15],Z[4][15],Z[3][15],Z[2][15],Z[1][15],Z[0][15]},opcode);
	mux_8_1 m_16(Y[16],{Z[7][16],Z[6][16],Z[5][16],Z[4][16],Z[3][16],Z[2][16],Z[1][16],Z[0][16]},opcode);
	mux_8_1 m_17(Y[17],{Z[7][17],Z[6][17],Z[5][17],Z[4][17],Z[3][17],Z[2][17],Z[1][17],Z[0][17]},opcode);
	mux_8_1 m_18(Y[18],{Z[7][18],Z[6][18],Z[5][18],Z[4][18],Z[3][18],Z[2][18],Z[1][18],Z[0][18]},opcode);
	mux_8_1 m_19(Y[19],{Z[7][19],Z[6][19],Z[5][19],Z[4][19],Z[3][19],Z[2][19],Z[1][19],Z[0][19]},opcode);
	mux_8_1 m_20(Y[20],{Z[7][20],Z[6][20],Z[5][20],Z[4][20],Z[3][20],Z[2][20],Z[1][20],Z[0][20]},opcode);
	mux_8_1 m_21(Y[21],{Z[7][21],Z[6][21],Z[5][21],Z[4][21],Z[3][21],Z[2][21],Z[1][21],Z[0][21]},opcode);
	mux_8_1 m_22(Y[22],{Z[7][22],Z[6][22],Z[5][22],Z[4][22],Z[3][22],Z[2][22],Z[1][22],Z[0][22]},opcode);
	mux_8_1 m_23(Y[23],{Z[7][23],Z[6][23],Z[5][23],Z[4][23],Z[3][23],Z[2][23],Z[1][23],Z[0][23]},opcode);
	mux_8_1 m_24(Y[24],{Z[7][24],Z[6][24],Z[5][24],Z[4][24],Z[3][24],Z[2][24],Z[1][24],Z[0][24]},opcode);
	mux_8_1 m_25(Y[25],{Z[7][25],Z[6][25],Z[5][25],Z[4][25],Z[3][25],Z[2][25],Z[1][25],Z[0][25]},opcode);
	mux_8_1 m_26(Y[26],{Z[7][26],Z[6][26],Z[5][26],Z[4][26],Z[3][26],Z[2][26],Z[1][26],Z[0][26]},opcode);
	mux_8_1 m_27(Y[27],{Z[7][27],Z[6][27],Z[5][27],Z[4][27],Z[3][27],Z[2][27],Z[1][27],Z[0][27]},opcode);
	mux_8_1 m_28(Y[28],{Z[7][28],Z[6][28],Z[5][28],Z[4][28],Z[3][28],Z[2][28],Z[1][28],Z[0][28]},opcode);
	mux_8_1 m_29(Y[29],{Z[7][29],Z[6][29],Z[5][29],Z[4][29],Z[3][29],Z[2][29],Z[1][29],Z[0][29]},opcode);
	mux_8_1 m_30(Y[30],{Z[7][30],Z[6][30],Z[5][30],Z[4][30],Z[3][30],Z[2][30],Z[1][30],Z[0][30]},opcode);
	mux_8_1 m_31(Y[31],{Z[7][31],Z[6][31],Z[5][31],Z[4][31],Z[3][31],Z[2][31],Z[1][31],Z[0][31]},opcode);

endmodule
