`include "multiplexers.v"

/* 64 bit Barrel Shifter using 64:1 Multiplexer*/
module barrelShift_64(Y, X, D);

	// I/O Port Declarations
	output[63:0] Y;
	input[63:0] X;
	input[5:0] D;

	// row of multiplexers
	mux_64_1 m64_0(Y[63], {X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63]}, D);
	mux_64_1 m64_1(Y[62], {X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62]}, D);
	mux_64_1 m64_2(Y[61], {X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61]}, D);
	mux_64_1 m64_3(Y[60], {X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60]}, D);
	mux_64_1 m64_4(Y[59], {X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59]}, D);
	mux_64_1 m64_5(Y[58], {X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58]}, D);
	mux_64_1 m64_6(Y[57], {X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57]}, D);
	mux_64_1 m64_7(Y[56], {X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56]}, D);
	mux_64_1 m64_8(Y[55], {X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55]}, D);
	mux_64_1 m64_9(Y[54], {X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54]}, D);
	mux_64_1 m64_10(Y[53], {X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53]}, D);
	mux_64_1 m64_11(Y[52], {X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52]}, D);
	mux_64_1 m64_12(Y[51], {X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51]}, D);
	mux_64_1 m64_13(Y[50], {X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50]}, D);
	mux_64_1 m64_14(Y[49], {X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49]}, D);
	mux_64_1 m64_15(Y[48], {X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48]}, D);
	mux_64_1 m64_16(Y[47], {X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47]}, D);
	mux_64_1 m64_17(Y[46], {X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46]}, D);
	mux_64_1 m64_18(Y[45], {X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45]}, D);
	mux_64_1 m64_19(Y[44], {X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44]}, D);
	mux_64_1 m64_20(Y[43], {X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43]}, D);
	mux_64_1 m64_21(Y[42], {X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42]}, D);
	mux_64_1 m64_22(Y[41], {X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41]}, D);
	mux_64_1 m64_23(Y[40], {X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40]}, D);
	mux_64_1 m64_24(Y[39], {X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39]}, D);
	mux_64_1 m64_25(Y[38], {X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38]}, D);
	mux_64_1 m64_26(Y[37], {X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37]}, D);
	mux_64_1 m64_27(Y[36], {X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36]}, D);
	mux_64_1 m64_28(Y[35], {X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35]}, D);
	mux_64_1 m64_29(Y[34], {X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34]}, D);
	mux_64_1 m64_30(Y[33], {X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33]}, D);
	mux_64_1 m64_31(Y[32], {X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32]}, D);
	mux_64_1 m64_32(Y[31], {X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31]}, D);
	mux_64_1 m64_33(Y[30], {X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30]}, D);
	mux_64_1 m64_34(Y[29], {X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29]}, D);
	mux_64_1 m64_35(Y[28], {X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28]}, D);
	mux_64_1 m64_36(Y[27], {X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27]}, D);
	mux_64_1 m64_37(Y[26], {X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26]}, D);
	mux_64_1 m64_38(Y[25], {X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25]}, D);
	mux_64_1 m64_39(Y[24], {X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24]}, D);
	mux_64_1 m64_40(Y[23], {X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23]}, D);
	mux_64_1 m64_41(Y[22], {X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22]}, D);
	mux_64_1 m64_42(Y[21], {X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21]}, D);
	mux_64_1 m64_43(Y[20], {X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20]}, D);
	mux_64_1 m64_44(Y[19], {X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19]}, D);
	mux_64_1 m64_45(Y[18], {X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18]}, D);
	mux_64_1 m64_46(Y[17], {X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17]}, D);
	mux_64_1 m64_47(Y[16], {X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16]}, D);
	mux_64_1 m64_48(Y[15], {X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15]}, D);
	mux_64_1 m64_49(Y[14], {X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14]}, D);
	mux_64_1 m64_50(Y[13], {X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13]}, D);
	mux_64_1 m64_51(Y[12], {X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12]}, D);
	mux_64_1 m64_52(Y[11], {X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11]}, D);
	mux_64_1 m64_53(Y[10], {X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10]}, D);
	mux_64_1 m64_54(Y[9], {X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9]}, D);
	mux_64_1 m64_55(Y[8], {X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8]}, D);
	mux_64_1 m64_56(Y[7], {X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6],X[7]}, D);
	mux_64_1 m64_57(Y[6], {X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5],X[6]}, D);
	mux_64_1 m64_58(Y[5], {X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4],X[5]}, D);
	mux_64_1 m64_59(Y[4], {X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3],X[4]}, D);
	mux_64_1 m64_60(Y[3], {X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2],X[3]}, D);
	mux_64_1 m64_61(Y[2], {X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1],X[2]}, D);
	mux_64_1 m64_62(Y[1], {X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0],X[1]}, D);
	mux_64_1 m64_63(Y[0], {X[1],X[2],X[3],X[4],X[5],X[6],X[7],X[8],X[9],X[10],X[11],X[12],X[13],X[14],X[15],X[16],X[17],X[18],X[19],X[20],X[21],X[22],X[23],X[24],X[25],X[26],X[27],X[28],X[29],X[30],X[31],X[32],X[33],X[34],X[35],X[36],X[37],X[38],X[39],X[40],X[41],X[42],X[43],X[44],X[45],X[46],X[47],X[48],X[49],X[50],X[51],X[52],X[53],X[54],X[55],X[56],X[57],X[58],X[59],X[60],X[61],X[62],X[63],X[0]}, D);

endmodule