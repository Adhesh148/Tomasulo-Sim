`include "fpAdd.v"

module top;
	reg[31:0] X1,X2;
	wire[31:0] X3;

	fpADD_32 fp_0 (X3 ,X1, X2);

	// Setup the monitoring for the signal values
	initial
	begin
		$monitor($time," X1 = %b,  X2 = %b --- X3 = %b\n",X1,X2,X3);
		$dumpfile("fpa.vcd");
		$dumpvars;
	end

	// Simulate the inputs
	initial
	begin
		X1 = 0; X2 = 0;

		#5 X1 = 32'b01000000010001100110011001100110; X2 = 32'b01000000111000000000000000000000;

		// 9.75 + 0.5625 = 10.3125
		#5 X2 = 32'b01000001000111000000000000000000; X1 = 32'b00111111000100000000000000000000;

		// 4 + 0.1  = 4.09999990463
		#5 X2 = 32'b01000000100000000000000000000000; X1 = 32'b00111101110011001100110011001101;

		// 4 - 0.25 = 3.75
		#5 X1 = 32'b01000000100000000000000000000000; X2 = 32'b10111110100000000000000000000000;

		// 4.13000011444 + 2.40000009537 = 6.53000020981
		#5 X1 = 32'b01000000100001000010100011110110; X2 = 32'b01000000000110011001100110011010;

		// -4 + 0.25 = -3.75
		#5 X1 = 32'b11000000100000000000000000000000; X2 = 32'b00111110100000000000000000000000;

		// 4 - 6.25 = -2.25
		#5 X1 = 32'b01000000100000000000000000000000; X2 = 32'b11000000110010000000000000000000;

		// 4 - 4 = 0
		#5 X1 = 32'b01000000100000000000000000000000; X2 = 32'b11000000100000000000000000000000;

		// -4 + (-4.0078125)
		#5 X1 = 32'b11000000100000000000000000000000; X2 = 32'b11000000100000000100000000000000;

		// -2312.12 + (-142.912)
		#5 X1 = 32'b11000101000100001000000111101100; X2 = 32'b11000011000011101110100101111001;
		
		// -990.99 + 0.99
		#5 X1 = 32'b11000100011101111011111101011100; X2 = 32'b00111111011111010111000010100100;

		//  inf  + 3
		#5 X1 = 32'b01111111100000000000000000000000; X2 = 32'b01000000010000000000000000000000;

		// 7.37869762948e+19 + 4.42721857769e+20 = 5.16508834064e+20
		#5 X1 = 32'b01100000100000000000000000000000; X2 = 32'b01100001110000000000000000000000;

		// 7.37869762948e+19 - 4.42721857769e+20 = -3.68934881474e+20
		#5 X1 = 32'b01100000100000000000000000000000; X2 = 32'b11100001110000000000000000000000;

		//  inf  + inf = inf
		#5 X1 = 32'b01111111100000000000000000000000; X2 = 32'b01111111100000000000000000000000;

	end

endmodule